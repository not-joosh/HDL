/*********************************************************
*	File: 				tb_4-BitAdder.v
*	Author: 				Josh Ratificar
*	Class:				CpE 3101L Introduction to HDL
*	Group/Schedule:	Friday, 7:30 AM to 10:30 AM
*	Description:		Testbench file for 4-BitAdder.v
*********************************************************/
`timescale 1 ns/ 1 ps
module tb_FourBitAdder();
	// all inputs to UUT are declared as reg type 
	reg		[3:0] A, B;
	reg		C_in;
	wire		[3:0] S;
	wire		C_out;
	// instantiate UUT with implicit oprt mapping
	FourBitAdder UUT (A[3:0], B[3:0], C_in, S[3:0], C_out);
	
	// generate stimuli
	initial
	begin
		A =  4'd0;	B = 4'd0;	C_in = 0;	#10
		A =  4'd3;	B = 4'd8;	C_in = 1;	#10
		A =  4'd11;	B = 4'd3;	C_in = 0;	#10
		A =  4'd12;	B = 4'd6;	C_in = 0;	#10
		A =  4'd5;	B = 4'd4;	C_in = 1;	#10
		A =  4'd1;	B = 4'd9;	C_in = 0;	#10
		A =  4'd15;	B = 4'd15;	C_in = 0;	#10
		A =  4'd15;	B = 4'd15;	C_in = 1;	#10
		$stop;
	end
endmodule
